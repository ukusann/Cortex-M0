`timescale 1ns / 1ps


module ControlUnit(
    input wire clk,
    input wire rst

    );
endmodule
